library verilog;
use verilog.vl_types.all;
entity sisc_tb_2 is
    generic(
        tclk            : real    := 10.000000
    );
end sisc_tb_2;
